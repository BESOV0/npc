module ysyx_22050598_IFU(
input clk,
input rst,
input [63:0] pc,
output [31:0] pc_inst,
//output next_pc
);

 
 







endmodule
